/* Using two 8x1 mux and 2x1 mux */

module mux_16x1(out, i, s);

input [15:0] i;
input [3:0] s;

output out;

/* Using 8x1 and 2x1
wire out1, out2;

mux_8x1 m1(out1, i[7:0], s[2:0]);
mux_8x1 m2(out2, i[15:8], s[2:0]);

mux_2x1 m3(out, out1, out2, s[3]);

*/

/* Using 4x1 mux */

wire [3:0] w;

mux_4x1 mux1(w[0], i[3:0], s[1:0]);
mux_4x1 mux2(w[1], i[7:4], s[1:0]);
mux_4x1 mux3(w[2], i[11:8], s[1:0]);
mux_4x1 mux4(w[3], i[15:12], s[1:0]);

mux_4x1 mux5(out, w, s[3:2]);

endmodule


/*
module testbench;

reg [15:0] i;
reg [3:0] s;

wire out;

mux_16x1 m1(out, i, s);

initial begin

     s = 4'b0000; i = 16'b0000000000000001;
#100 s = 4'b0001; i = 16'b0000000000000010;
#100 s = 4'b0010; i = 16'b0000000000000100;
#100 s = 4'b0011; i = 16'b0000000000001000;
#100 s = 4'b0100; i = 16'b0000000000010000;
#100 s = 4'b0101; i = 16'b0000000000100000;
#100 s = 4'b0110; i = 16'b0000000001000000;
#100 s = 4'b0111; i = 16'b0000000010000000;
#100 s = 4'b1000; i = 16'b0000000100000000;
#100 s = 4'b1001; i = 16'b0000001000000000;
#100 s = 4'b1010; i = 16'b0000010000000000;
#100 s = 4'b1011; i = 16'b0000100000000000;
#100 s = 4'b1100; i = 16'b0001000000000000;
#100 s = 4'b1101; i = 16'b0010000000000000;
#100 s = 4'b1110; i = 16'b0100000000000000;
#100 s = 4'b1111; i = 16'b1000000000000000;

end

endmodule
*/