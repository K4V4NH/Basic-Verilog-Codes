module aoitb;
reg a1,a2,b1,b2;
wire o;
Aoi go(a1,a2,b1,b2,o);
initial begin
{a1,a2,b1,b2} =4'b0000;
#100 {a1,a2,b1,b2} =4'b0001;
#100 {a1,a2,b1,b2} =4'b0010;
#100 {a1,a2,b1,b2} =4'b0011;
#100 {a1,a2,b1,b2} =4'b0100;
#100 {a1,a2,b1,b2} =4'b0101;
#100 {a1,a2,b1,b2} =4'b0110;
#100 {a1,a2,b1,b2} =4'b0111;
#100 {a1,a2,b1,b2} =4'b1000;
#100 {a1,a2,b1,b2} =4'b1001;
#100 {a1,a2,b1,b2} =4'b1010;
#100 {a1,a2,b1,b2} =4'b1011;
#100 {a1,a2,b1,b2} =4'b1100;
#100 {a1,a2,b1,b2} =4'b1101;
#100 {a1,a2,b1,b2} =4'b1110;
#100 {a1,a2,b1,b2} =4'b1111;
end
endmodule
 